`timescale 1ns/1ps

module APB_SLAVE(PCLK, PRESETn, PADDR, PSELx, PENABLE, PWRITE, PWDATA, PREADY, PSLVERR, PRDATA);
parameter DW = 32;
parameter AW = 32;
parameter DELAY =2;

input PCLK, PRESETn, PSELx, PENABLE, PWRITE;
input [AW-1:0] PADDR;
input [DW-1:0] PWDATA;
output PREADY, PSLVERR;
output [DW-1:0] PRDATA;

wire [DW-1:0] WDATA, RDATA;
wire [AW/2-1:0] ADDR;
wire 			W_ENABLE;


//APB_SLAVE_Mealy   slave(PCLK, PRESETn, PADDR, PSELx, PENABLE, PWRITE, PWDATA, PREADY, PSLVERR, ADDR, W_ENABLE, pWDATA);
APB_SLAVE_Mealy   slave(PCLK, PRESETn, PADDR, PSELx, PENABLE, RDATA, PWRITE, PRDATA, PWDATA, PREADY, PSLVERR, ADDR, W_ENABLE, WDATA);
Reg_File 		register(PCLK, W_ENABLE, PRESETn, ADDR, WDATA, RDATA);


endmodule